
`define LENGTH 16